/afs/ee.cooper.edu/user/d/david.yang/VLSI_tsmc65/yangd_lvs/netlist